* 134-158MHz Chebychev bandpass filter, simulated from:
* https://markimicrowave.com/technical-resources/tools/lc-filter-design-tool/
* 3rd order, conventional shunt first, 134 low cutoff, 158 high
* cutoff, .10db ripple in passband, 50 ohm input, 50 ohm output
* impedance.  input | output | | .SUBCKT Filt144MHz in out

*                  input
*                  |   output
*                  |   |
.SUBCKT Filt144MHz in  out

* Comments above are the exact values from the filter tool.
* Value used are available inductors and capacitors.

* 136.8p
C1	in  0   136p
* 8.745n
L1	in  0   8.7n

* 3.145p
C2	in  a1 3.1p
* 380.4
L2	a1  out 380n

C3	out 0   136p
L3	out 0   8.7n

* Avoid issues with series inductors, they result in:
* Warning: singular matrix:  check node l.x1.l4b#branch
* Warning: True gmin stepping failed
* This add a series resistor on all inductors.
.option rseries = 1.0e-4

.ENDS

V1 0 in dc 0 AC 1 sin(0 1 146MEG 0 0 0)
Rsrc in in1 50

X1 in1 out Filt144MHz

Rload out 0 50

.control
*tran 1ns 102000ns 101000ns
*plot v(in1), v(out)
ac lin 50000 120Meg 180Meg
plot db((vm(out)^2/50)/(vm(in1) * i(v1)))
.endc

.end
