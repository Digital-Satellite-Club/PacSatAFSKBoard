* 123-173MHz Chebychev bandpass filter, simulated from:
* https://markimicrowave.com/technical-resources/tools/lc-filter-design-tool/
* 3rd order, conventional shunt first, 123 low cutoff, 173 high
* cutoff, .10db ripple in passband, 50 ohm input, 50 ohm output
* impedance.

*                  input
*                  |   output
*                  |   |
.SUBCKT Filt144MHz in  out

* Comments above are the exact values from the filter tool.
* Value used are available inductors and capacitors.

* 65.57p
C1	in  0   68p
* 18.13n
L1	in  b1  18n
R1      b1  0   .078

* 6.519p
C2	in  a1  6.5p
* 182.6
L2	a1  a2  180n
R2	a2  b3  .64

C3	b3  0   68p
L3	b3  b2   18n
R3      b2  0   .078

* Impedance matching network
L4      b3  b4  91n
R4      b4  out .576
C4      out 0   6.5p

.ENDS

V1 0 in dc 0 AC 1 sin(0 1 146MEG 0 0 0)
Rsrc in in1 50

X1 in1 out Filt144MHz

Cload out out1 13.6p

* Used for current measurement.
Vload out1 out2 DC 0 AC 0

* Input impedance of the LNA
Rload out2 0 142.4

.control
*tran 1ns 102000ns 101000ns
*plot v(in1), v(out)
ac lin 50000 100Meg 500Meg
plot db((v(out1) * i(Vload)) / (vm(in1) * i(V1)))
.endc

.end
