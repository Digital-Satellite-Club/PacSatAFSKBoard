* 460MHz Elliptic lowpass filter, simulated from:
* https://markimicrowave.com/technical-resources/tools/lc-filter-design-tool/
* 5rd order, shunt first, 460MHz cutoff, .10db ripple in passband, 50
* ohm input, 50 ohm output impedance, 50dB stopband attenuation.

*                     input
*                     |   output
*                     |   |
.SUBCKT ImpMatchPAOut in  out

* Impedance matching network
*Lin     in   inx  10.9n
*Rin     inx  out  .078
*Cout    out  0    19.5p

* The above are the calculated values.  For some reason they don't
* work well in simulation.  The below work much better in simulation.
* I need to figure out why.

Lin     in   inx  .2n
Rin     inx  out  .078
Cout    out  0    3.5p

.ENDS

*                  input
*                  |   output
*                  |   |
.SUBCKT Filt440MHz in  out

* 7.32p
C1	in   0   7.32p

* 21.71n
L2	in  a1  21.71n
R2      a1  a2   .078
* 767.6f
C2	in  a2  .768p

* 11.84p
C3	a2  0   11.84p

* 17.96n
L4	a2  a3  17.96n
R4	a3  out .078
* 2.16p
C4	a2  out 2.16p

* 6.2p
C5	out 0   6.2p

.ENDS

V1 0 ina dc 0 AC 1 sin(0 1 435MEG 0 0 0)

Rsrc ina ina1  6.23
Csrc ina1 in 27p
*Rsrc ina in  50

X1 in  im1 ImpMatchPAOut

* Used for current measurement.
Vm1 im1 im2 AC 0 DC 0

X2 im2 out Filt440MHz

* Used for current measurement.
Vmout out out2 DC 0 AC 0

Rload out2 0    50
*Rload out2 out1 6.23
*Cload out1 0    27p

.control
*tran 1ns 102000ns 101000ns
*plot v(in1), v(out)

ac lin 5000 400Meg 470Meg
plot vr(out) vi(out) vp(out)

ac lin 50000 300Meg 1000Meg
plot db((v(out) * i(Vmout)) / (vm(in) * i(V1)))
plot db((v(im1) * i(Vm1)) / (vm(in) * i(V1)))
*plot db((v(out) * i(Vmout)) / (vm(im1) * i(Vm1)))

*plot db(v(out) * i(Vload)) db(v(in2) * i(VLoad1)) db(vm(in1) * i(V1))
.endc

.end
