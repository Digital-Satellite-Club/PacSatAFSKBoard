* RF input filter from the antenna to the LNA

* Unless otherwise mentioned, assume all inductors have a Q of around 35
* at 144MHz.  This is a pretty good assumption for the Coilcraft 0603DC
* inductors.

*                  input
*                  |   output
*                  |   |
.SUBCKT Filt144MHz in  out

* Comments above are the exact values from the filter tool.
* Value used are available inductors and capacitors.

.if (1)
* 176MHz Elliptic lowpass filter, shunt first, with 50dB stopband
* attenuation and 1dB ripple in the passband.  50ohm input and output.

* This is the inductor used to bleed off static from the antenna
L0	in	b0	470n
R0	b0	0	10k

* 35.62
C1	in	0	36p

* 1.203p
C2	in	out	1p
* 43.03n
L1	in	b1	43n
Rl1	b1	out	1.15
Cl1	in	out	.18p

C3	out	0	36p

.endif

.if (0)
* 123-173MHz Chebychev bandpass filter, simulated from:
* https://markimicrowave.com/technical-resources/tools/lc-filter-design-tool/
* 3rd order, conventional shunt first, 123MHz low cutoff, 173MHz high
* cutoff, .10db ripple in passband, 50 ohm input, 50 ohm output
* impedance.

* 65.57p
C1	in	0	68p
* 18.13n
L1	in	b1	18n
R1      b1	0	.5

* 6.519p
C2	in	a1	6.5p
* 182.6 * Coilcraft 0805CS series has a Q of around 50
L2	a1	a2	180n
R2	a2	out	3.39

C3	out	0	68p
L3	out	b2	18n
R3      b2	0	.5
.endif

.ENDS

.SUBCKT ImpMatchLNAIn in out

* TX LNA input matcher
L1	in	a1	91n
* Coilcraft 0805CS series has a Q of around 50
Rl1	a1	out	1.7
Cl1	in	out	.16p
C1	out	0	6.5p

.ENDS


V1 0 in dc 0 AC 1 sin(0 1 146MEG 0 0 0)
Rsrc in in1 50

X1 in1 im1 Filt144MHz

X2 im1 out ImpMatchLNAin

Cload out out1 13.6p

* Used for current measurement.
Vload out1 out2 DC 0 AC 0

* Input impedance of the LNA
Rload out2 0 142.4

.control
*tran 1ns 102000ns 101000ns
*plot v(in1), v(out)
ac lin 50000 1Meg 500Meg
plot db((v(out1) * i(Vload)) / (vm(in1) * i(V1)))
.endc

.end
