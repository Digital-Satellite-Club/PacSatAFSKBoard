* 460MHz Elliptic lowpass filter, simulated from:
* https://markimicrowave.com/technical-resources/tools/lc-filter-design-tool/
* 5rd order, shunt first, 460MHz cutoff, .10db ripple in passband, 50
* ohm input, 50 ohm output impedance, 50dB stopband attenuation.

*                     input
*                     |   output
*                     |   |
.SUBCKT ImpMatchPAOut in  out

* Impedance matching network
C1     in     out 110p
L1     inx    a3  6.9n
R1     a3     0   .078

.ENDS

*                  input
*                  |   output
*                  |   |
.SUBCKT Filt440MHz in  out

* 7.32p
C1	in   0   7.3p

* 21.71n
L2	in  a1  22n
R2      a1  a2  .078
* 767.6f
C2	in  a2  .75p

* 11.84p
C3	a2  0   12p

* 17.96n
L4	a2  a3  18n
R4	a3  out .078
* 2.16p
C4	a2  out 2.2p

* 6.2p
C5	out 0   6.2p

.ENDS

V1 ina 0 dc 0 AC 1 sin(0 1 435MEG 0 0 0)

Rsrc ina  ina1 6.23
Csrc ina1 ina2 27p
*Rsrc ina ina1  50

* Used for current measurement.
Vmin ina2 in AC 0 DC 0

X1 in  im1 ImpMatchPAOut


* Used for current measurement.
Vm1 im1 im2 AC 0 DC 0

X2 im2 out Filt440MHz

* Used for current measurement.
Vmout out out2 DC 0 AC 0

Rload out2 0    50
*Rload out2 out1 6.23
*Cload out1 0    27p

.control
*tran 1ns 102000ns 101000ns
*plot v(in1), v(out)

ac lin 50000 3Meg 1000Meg
plot db((v(out) * i(Vmout)) / (vm(ina1) * i(V1)))
plot vr(out) vi(out) vp(out)

.endc

.end
