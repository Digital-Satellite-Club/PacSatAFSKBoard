* 140-150MHz Elliptic bandpass filter, simulated from:
* https://markimicrowave.com/technical-resources/tools/lc-filter-design-tool/
* 3rd order, conventional shunt first, 140 low cutoff, 150 high
* cutoff, .10db ripple in passband, 50 ohm input, 50 ohm output
* impedance, 50.42dB stopband attenuation

* Realization with real components brings about 2.5dB loss and shifts
* the frequency to 140-152MHz 3dB points.

.SUBCKT ImpMatchLNAOut in out

* TX LNA output matcher
C1   in     0       11p
L1   in     a1      47n
R1   a1     out     .2

.ENDS

*                    input
*                    |   output
*                    |   |
.SUBCKT FiltEl144MHz in  out

* Comments above are the exact values from the filter tool.
* Value used are available inductors and capacitors.

* Note that almost all of the loss is in R1 and R4.  R2 and R3 make
* very little contribution to the loss.  If inductors could be found
* that have lower series resistance it would greatly improve the loss
* in the filter.  Using two larger inductors in parallel results in
* lowering the series resistance from 46m to 26.5m, making about 2dB
* improvement.

.if (1)
* 322.4p
C1	in	0	320p
* 3.742n * 2% Q=68 0402DC-3N7XGRW
*L1	in	b1	3.7n
*R1	b1	0	.046
* 7.5n 2% Q=88 0603DC-7N5XGRW
L1a	in	b1a	7.5n
R1a	b1a	0	.053
L1b	in	b1b	7.5n
R1b	b1b	0	.053

* 13.25p
C2	in	a1	13p
* 60.45n * 62n 2% Q=70 LQW2BAN62NG00L 0805
L2	in	a2	62n
R2	a2	a1	.120

* 19.95p
C3	a1	out	20p
* 91.06n * 91n 2% Q=70 LQW2BAN91NG00L 0805
L3	a1	a4	91n
R3	a4	out	.210

* Same as first values above.
C4	out	0	320p
*L4	out	b2	3.7n
*R4	b2	0	.046
L4a	out	b2a	7.5n
R4a	b2a	0	.053
L4b	out	b2b	7.5n
R4b	b2b	0	.053
.endif

.if (0)
* This is a 3rd order Chebychev bandpass filter direct coupled, shunt
* capacitor, 140 to 150MHz .1dB ripple in the passband, 50 ohms input
* and output impedance.  The direct coupled inductor is 91nH.
*
* This has slightly less loss than the Elliptic filter, but not as
* good performance.  The nice thing is you pick a single inductor
* value, so dealing with the inductor isn't so hard.  Performance
* is more important than loss at this point.

* 
C1	in	0	62.13p
*
C2	in	a1	17.69p
* 
L1	a1	a2	91n
R1	a2	a3	.210
*
C3	a3	0	208.7p
*
C4	a3	a4	15.14p
*
L2	a4	a5	91n
R2	a5	a6	.210
*
C5	a6	0	208.7p
*
C6	a6	a7	17.69p
* 
L3	a7	a8	91n
R3	a8	out	.210
*
C7	out	0	62.13p
.endif

.ENDS

V1 in 0 dc 0 AC 1 sin(0 1 146MEG 0 0 0)

* LNA output impedance and measurement voltage source
Rsrc in     in0  86.6
* Used for current measurement
Vm1  in0  in1  DC 0 AC 0
* -1.88 ohms at 145MHz
Csrc in1    in2  583p

X1 in2 im1 ImpMatchLNAOut

Vm2  im1  im2  DC 0 AC 0

X2 im2 out FiltEl144MHz

* Used for current measurement.
Vload out out2 DC 0 AC 0

* Input impedance of the LNA
Rload out2 0   50

.control
*tran 1ns 102000ns 101000ns
*plot v(in1), v(out)
ac lin 50000 100Meg 200Meg
plot db((v(out) * i(Vload)) / (v(in0) * i(Vm1)))
.endc

.end
