*
* This contains small simulations of the iput and output impedance
* matching circuits in the LNA and PA sections.  Modify the if
* statements to get the one you want, make sure to look at the
* graph with the right frequencies!
*
* Also remember that on the output side, the load side of the match
* is looking into the PA/LNA device.  So it's backwards.
*

*.option rseries = 1.0e-4

.param pa_in=0

.SUBCKT ImpMatchPAIn in vmin1 vmin2 vmout1 vmout2

Rsrc in     vmin1  50

* TX PA input matcher
C1   vmin2  0      39p
L1   vmin2  a1a    18n
R1   a1a    a1     .078

* -37.7 ohms at 435MHz
Cout a1     vmout1 9.6p
Rout vmout2 0      1.87

.ENDS

.SUBCKT ImpMatchPAOut in vmin1 vmin2 vmout1 vmout2

Rsrc in     vmin1  6.23
* -13.3 ohms at 435MHz
Csrc vmin2  a1     27.5p

* Set the DC bias between two capacitors.
Rb1  a1     0      1Meg

* Impedance matching network
* TX PA output matcher
C1   a1     vmout1 110p
L1   vmout1 a3     6.9n
R1   a3     0      .063

Rout vmout2 0      50

.ENDS

.SUBCKT ImpMatchLNAIn in vmin1 vmin2 vmout1 vmout2

Rsrc in     vmin1  50

* TX LNA input matcher
L1   vmin2  a2   91n
R1   a2     a1   2.45
C1   a1     0    6.5p

* -80.8 ohms at 145MHz
Cout a1     vmout1 13.6p
Rout vmout2 0      142.4

.ENDS

.SUBCKT ImpMatchLNAOut in vmin1 vmin2 vmout1 vmout2

Rsrc in     vmin1  86.6
* -1.88 ohms at 145MHz
Csrc vmin2  a1     583p

* Set the DC bias between two capacitors.
Rb1  a1     0      1Meg

* TX LNA output matcher
C1   a1     0       11p
L1   a1     a2      47n
R1   a2     vmout1  .2

Rout vmout2 0      50

.ENDS

.param m = 0

.if (m == 1)
X1 in vmin1 vmin2 vmout1 vmout2 ImpMatchPAIn
.endif
.if (m == 2)
X1 in vmin1 vmin2 vmout1 vmout2 ImpMatchPAOut
.endif
.if (m == 3)
X1 in vmin1 vmin2 vmout1 vmout2 ImpMatchLNAIn
.endif
.if (m == 4)
X1 in vmin1 vmin2 vmout1 vmout2 ImpMatchLNAOut
.endif

V1 in 0 dc 0 AC 1 sin(1 0 435MEG 0 0 0)

* For current measurement
Vmin  vmin1  vmin2  dc 0 ac 0

* For current measurement
Vmout vmout1 vmout2 dc 0 ac 0

.control

alterparam m = 1
reset
ac lin 5000 1Meg 1000meg
plot title "PA Input" db((v(vmout1) * i(Vmout)) / (v(vmin1) * i(Vmin)))
plot title "PA Input" vi(vmin1)

alterparam m = 2
reset
ac lin 5000 1Meg 1000meg
plot title "PA Output" db((v(vmout1) * i(Vmout)) / (v(vmin1) * i(Vmin)))
plot title "PA Output" vi(vmin1)

alterparam m = 3
reset
ac lin 5000 1Meg 400meg
plot title "LNA Input" db((v(vmout1) * i(Vmout)) / (v(vmin1) * i(Vmin)))
plot title "LNA Input" vi(vmin1)

alterparam m = 4
reset
ac lin 5000 1Meg 400meg
plot title "LNA Output" db((v(vmout1) * i(Vmout)) / (v(vmin1) * i(Vmin)))
plot title "LNA Output" vi(vmin1)

.endc

.end
